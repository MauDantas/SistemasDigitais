module calculadoraBCD(A,B,d,u,o1,o0,sinal);
	input [2:0]A,B;
	input o1,o0;
	wire [6:0]F;
	output[3:0]d,u;
	output sinal;
	
	calculadora calculadora(A,B,F,o1,o0);
	
	assign u =F[6]?(F[3:0]*(-1)):(((F[5]&&F[4])||(F[5:1]== 5'b10011)||(F[5:1]== 5'b01110)||(F[5:1]== 5'b01001)||(F[5:1]== 5'b00100))?(4'b1000+F[0]):(((F[5:1]== 5'b10111)||(F[5:1]== 5'b10010)||(F[5:1]== 5'b01101)||(F[5:1]== 5'b01000)||(F[5:1]== 5'b00011))?(4'b0110+F[0]):(((F[5:1]== 5'b10110)||(F[5:1]== 5'b10001)||(F[5:1]== 5'b01100)||(F[5:1]== 5'b00111)||(F[5:1]== 5'b00010))?(4'b0100+F[0]):(((F[5:1]== 5'b10101)||(F[5:1]== 5'b10000)||(F[5:1]== 5'b01011)||(F[5:1]== 5'b00110)||(F[5:1]== 5'b00001))?(4'b0010+F[0]):(4'b0000+F[0])))));
	assign d =F[6]?(4'b0000):(F[5]?(F[4]?(4'b0100):(F[3]?(4'b0100):(4'b011))):((&F[4:1])?(4'b0011):((F[3]&&F[4])?(4'b0010):((F[4]||(F[3]&&(F[2]||F[1])))?(4'b0001):(4'b0000)))));
	buf b1(sinal,F[6]);

endmodule
